`include "APB/apb_if.sv"
`include "APB/apb_pkt.sv"
`include "APB/apb_master_driver.sv"
`include "APB/apb_master_monitor.sv"
`include "APB/apb_master_seq.sv"
`include "APB/apb_master_sequencer.sv"
`include "APB/apb_master_config.sv"
`include "APB/apb_master_agent.sv"
