basava

